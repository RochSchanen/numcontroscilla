-- ########################################################

-- file: fpga_bench.vhd
-- content: bench to simulate fpga code
-- Created: 2024 july 28
-- Author: Roch Schanen
-- comments: simulate external clock, input and outputs ports.

-- ########################################################

-------------------------------------------------
--                FPGA BENCH
-------------------------------------------------

-- library IEEE;
-- use IEEE.STD_LOGIC_1164.ALL;

entity fpga_bench is

    -- ports

end fpga_bench;

architecture fpga_bench_arch of fpga_bench is

begin

    process
    begin

        -- nothing 
        report "done";
        wait;

    end process;

end fpga_bench_arch;

